LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM IS
    PORT
    (
        clk : IN std_logic;
        data_in : IN std_logic;
        reset : IN std_logic;
        student_id : OUT std_logic_vector(3 DOWNTO 0);
        current_state : OUT std_logic_vector(3 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE fsm OF FSM IS
    TYPE state_type IS (s0, s1, s2, s3, s4, s5, s6, s7, s8);
    SIGNAL yfsm : state_type;
BEGIN
    PROCESS (clk, reset)
    BEGIN
        IF reset = '1' THEN
            yfsm <= s0;
        ELSIF (clk'EVENT AND clk = '1') THEN
            CASE yfsm IS
                WHEN s0 =>
                    IF data_in = '0' THEN
                        yfsm <= s0;
                    ELSE
                        yfsm <= s1;
                    END IF;
                WHEN s1 =>
                    IF data_in = '0' THEN
                        yfsm <= s1;
                    ELSE
                        yfsm <= s2;
                    END IF;
                WHEN s2 =>
                    IF data_in = '0' THEN
                        yfsm <= s2;
                    ELSE
                        yfsm <= s3;
                    END IF;
                WHEN s3 =>
                    IF data_in = '0' THEN
                        yfsm <= s3;
                    ELSE
                        yfsm <= s4;
                    END IF;
                WHEN s4 =>
                    IF data_in = '0' THEN
                        yfsm <= s4;
                    ELSE
                        yfsm <= s5;
                    END IF;
                WHEN s5 =>
                    IF data_in = '0' THEN
                        yfsm <= s5;
                    ELSE
                        yfsm <= s6;
                    END IF;
                WHEN s6 =>
                    IF data_in = '0' THEN
                        yfsm <= s6;
                    ELSE
                        yfsm <= s7;
                    END IF;
                WHEN s7 =>
                    IF data_in = '0' THEN
                        yfsm <= s7;
                    ELSE
                        yfsm <= s8;
                    END IF;
                WHEN s8 =>
                    IF data_in = '0' THEN
                        yfsm <= s8;
                    ELSE
                        yfsm <= s0;
                    END IF;
            END CASE;
        END IF;
    END PROCESS;

    PROCESS (yfsm, data_in)
    BEGIN
        CASE yfsm IS
            WHEN s0 =>
                current_state <= "0000"; -- S0
                student_id <= "0101"; -- 5
            WHEN s1 =>
                current_state <= "0001"; -- S1
                student_id <= "0000"; -- 0
            WHEN s2 =>
                current_state <= "0010"; -- S2
                student_id <= "0001"; -- 1
            WHEN s3 =>
                current_state <= "0011"; -- S3
                student_id <= "0001"; -- 1
            WHEN s4 =>
                current_state <= "0100"; -- S4
                student_id <= "0101"; -- 5
            WHEN s5 =>
                current_state <= "0101"; -- S5
                student_id <= "1001"; -- 9
            WHEN s6 =>
                current_state <= "0110"; -- S6
                student_id <= "0100"; -- 4
            WHEN s7 =>
                current_state <= "0111"; -- S7
                student_id <= "0111"; -- 7
            WHEN s8 =>
                current_state <= "1000"; -- S8
                student_id <= "0010"; -- 2
        END CASE;
    END PROCESS;
END fsm;
